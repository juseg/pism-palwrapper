netcdf ccli { // Config overrides for Cordillera climate paper
variables:
        byte pism_overrides ;

    // Customized PDD parameters
                pism_overrides:pdd_factor_snow = 0.00304 ;
                pism_overrides:pdd_factor_snow_doc = "m K-1 day-1; measured on present glaciers in British Columbia by Shea et al 2009, J. Glac. 55 (189): 123-130" ;
                pism_overrides:pdd_factor_ice = 0.00459 ;
                pism_overrides:pdd_factor_ice_doc = "m K-1 day-1; measured on present glaciers in British Columbia by Shea et al 2009, J. Glac. 55 (189): 123-130" ;
                pism_overrides:pdd_std_dev = 3.068094 ;
                pism_overrides:pdd_std_dev_doc = "K; summer (JJA) average of monthly standard deviation over the entire domain computed from North American Regional Reanalysis data." ;
                pism_overrides:pdd_refreeze = 0.0 ;

    // Rebound model
                pism_overrides:bed_deformation_model = "lc" ;

    // Thickness calving
    pism_overrides:calving_methods = "thickness_calving" ;
    pism_overrides:thickness_calving_threshold = 200. ;
                pism_overrides:part_grid = "yes" ;
                pism_overrides:part_redist = "yes" ;

    // Constant geothermal heat flux
                pism_overrides:bootstrapping_geothermal_flux_value_no_var = 0.070 ;

    // SSA sliding
    pism_overrides:stress_balance_model = "ssa+sia" ;
                pism_overrides:till_effective_fraction_overburden = 0.05 ;
}
