netcdf pism_overrides {
variables:
        byte pism_overrides ;
                pism_overrides:calving_front_stress_boundary_condition = "yes" ;
                pism_overrides:calving_front_stress_boundary_condition_doc = "Apply CFBC condition as in [\\ref Albrechtetal2011, \\ref Winkelmannetal2010TCD].  May only apply to some stress balances; e.g. SSAFD as of May 2011.  If not set then a strength-extension is used, as in [\\ref BBssasliding]." ;
                pism_overrides:part_grid = "yes" ;
                pism_overrides:part_grid_doc = "apply partially filled grid cell scheme" ;
                pism_overrides:part_redist = "yes" ;
                pism_overrides:part_redist_doc = "for partially filled grid cell scheme, redistribute residuals Hresidual" ;
                pism_overrides:kill_icebergs = "yes" ;
                pism_overrides:kill_icebergs_doc = "identify and kill detached ice-shelf areas" ;
}
